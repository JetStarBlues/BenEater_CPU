library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.components_pk.all;


entity programMemoryXN is

	generic (

		X : integer
	);

	port (

		addr : in  std_logic_vector( N - 1 downto 0 );
		q    : out std_logic_vector( N - 1 downto 0 )
	);

end entity;


architecture ac of programMemoryXN is

	type rom_type is array( 0 to X - 1 ) of std_logic_vector( N - 1 downto 0 );
	
	constant rom : rom_type := (

		-- Increment ( OUT = OUT + 1 ) (datatype - uint8)
		--0 => "01010001",
		--1 => "01001111",
		--2 => "01010000",
		--3 => "00101111",
		--4 => "11100000",
		--5 => "01100011",

		-- Multiples of 3 ( OUT = 3x ) (datatype - uint8)
		--0 => "01010011",
		--1 => "01001111",
		--2 => "01010000",
		--3 => "00101111",
		--4 => "11100000",
		--5 => "01100011",

		-- Arithmetic test ( OUT = 5 + 2 - 15 ) (datatype - int8)
		--0  => "01010101",
		--1  => "01001111",
		--2  => "01010010",
		--3  => "01001110",
		--4  => "01011111",
		--5  => "01001101",
		--6  => "00011111",
		--7  => "00101110",
		--8  => "00111101",
		--9  => "11100000",
		--10 => "11110000",

		-- Hello world ( Greetings!\nIt's great to be awake!\n\n ) (datatype - ascii)
		  0 => "01011111",
		  1 => "01111111",
		  2 => "01111111",
		  3 => "01111111",
		  4 => "01111011",
		  5 => "11100000",
		  6 => "01011111",
		  7 => "01111111",
		  8 => "01111111",
		  9 => "01111111",
		 10 => "01111111",
		 11 => "01111111",
		 12 => "01111111",
		 13 => "01111001",
		 14 => "11100000",
		 15 => "01011111",
		 16 => "01111111",
		 17 => "01111111",
		 18 => "01111111",
		 19 => "01111111",
		 20 => "01111111",
		 21 => "01111011",
		 22 => "11100000",
		 23 => "01011111",
		 24 => "01111111",
		 25 => "01111111",
		 26 => "01111111",
		 27 => "01111111",
		 28 => "01111111",
		 29 => "01111011",
		 30 => "11100000",
		 31 => "01011111",
		 32 => "01111111",
		 33 => "01111111",
		 34 => "01111111",
		 35 => "01111111",
		 36 => "01111111",
		 37 => "01111111",
		 38 => "01111011",
		 39 => "11100000",
		 40 => "01011111",
		 41 => "01111111",
		 42 => "01111111",
		 43 => "01111111",
		 44 => "01111111",
		 45 => "01111111",
		 46 => "01111111",
		 47 => "01110000",
		 48 => "11100000",
		 49 => "01011111",
		 50 => "01111111",
		 51 => "01111111",
		 52 => "01111111",
		 53 => "01111111",
		 54 => "01111111",
		 55 => "01111111",
		 56 => "01110101",
		 57 => "11100000",
		 58 => "01011111",
		 59 => "01111111",
		 60 => "01111111",
		 61 => "01111111",
		 62 => "01111111",
		 63 => "01111111",
		 64 => "01111101",
		 65 => "11100000",
		 66 => "01011111",
		 67 => "01111111",
		 68 => "01111111",
		 69 => "01111111",
		 70 => "01111111",
		 71 => "01111111",
		 72 => "01111111",
		 73 => "01111010",
		 74 => "11100000",
		 75 => "01011111",
		 76 => "01111111",
		 77 => "01110011",
		 78 => "11100000",
		 79 => "01011010",
		 80 => "11100000",
		 81 => "01011111",
		 82 => "01111111",
		 83 => "01111111",
		 84 => "01111111",
		 85 => "01111101",
		 86 => "11100000",
		 87 => "01011111",
		 88 => "01111111",
		 89 => "01111111",
		 90 => "01111111",
		 91 => "01111111",
		 92 => "01111111",
		 93 => "01111111",
		 94 => "01111011",
		 95 => "11100000",
		 96 => "01011111",
		 97 => "01111111",
		 98 => "01111001",
		 99 => "11100000",
		100 => "01011111",
		101 => "01111111",
		102 => "01111111",
		103 => "01111111",
		104 => "01111111",
		105 => "01111111",
		106 => "01111111",
		107 => "01111010",
		108 => "11100000",
		109 => "01011111",
		110 => "01111111",
		111 => "01110010",
		112 => "11100000",
		113 => "01011111",
		114 => "01111111",
		115 => "01111111",
		116 => "01111111",
		117 => "01111111",
		118 => "01111111",
		119 => "01111101",
		120 => "11100000",
		121 => "01011111",
		122 => "01111111",
		123 => "01111111",
		124 => "01111111",
		125 => "01111111",
		126 => "01111111",
		127 => "01111111",
		128 => "01111001",
		129 => "11100000",
		130 => "01011111",
		131 => "01111111",
		132 => "01111111",
		133 => "01111111",
		134 => "01111111",
		135 => "01111111",
		136 => "01111011",
		137 => "11100000",
		138 => "01011111",
		139 => "01111111",
		140 => "01111111",
		141 => "01111111",
		142 => "01111111",
		143 => "01111111",
		144 => "01110111",
		145 => "11100000",
		146 => "01011111",
		147 => "01111111",
		148 => "01111111",
		149 => "01111111",
		150 => "01111111",
		151 => "01111111",
		152 => "01111111",
		153 => "01111011",
		154 => "11100000",
		155 => "01011111",
		156 => "01111111",
		157 => "01110010",
		158 => "11100000",
		159 => "01011111",
		160 => "01111111",
		161 => "01111111",
		162 => "01111111",
		163 => "01111111",
		164 => "01111111",
		165 => "01111111",
		166 => "01111011",
		167 => "11100000",
		168 => "01011111",
		169 => "01111111",
		170 => "01111111",
		171 => "01111111",
		172 => "01111111",
		173 => "01111111",
		174 => "01111111",
		175 => "01110110",
		176 => "11100000",
		177 => "01011111",
		178 => "01111111",
		179 => "01110010",
		180 => "11100000",
		181 => "01011111",
		182 => "01111111",
		183 => "01111111",
		184 => "01111111",
		185 => "01111111",
		186 => "01111111",
		187 => "01111000",
		188 => "11100000",
		189 => "01011111",
		190 => "01111111",
		191 => "01111111",
		192 => "01111111",
		193 => "01111111",
		194 => "01111111",
		195 => "01111011",
		196 => "11100000",
		197 => "01011111",
		198 => "01111111",
		199 => "01110010",
		200 => "11100000",
		201 => "01011111",
		202 => "01111111",
		203 => "01111111",
		204 => "01111111",
		205 => "01111111",
		206 => "01111111",
		207 => "01110111",
		208 => "11100000",
		209 => "01011111",
		210 => "01111111",
		211 => "01111111",
		212 => "01111111",
		213 => "01111111",
		214 => "01111111",
		215 => "01111111",
		216 => "01111110",
		217 => "11100000",
		218 => "01011111",
		219 => "01111111",
		220 => "01111111",
		221 => "01111111",
		222 => "01111111",
		223 => "01111111",
		224 => "01110111",
		225 => "11100000",
		226 => "01011111",
		227 => "01111111",
		228 => "01111111",
		229 => "01111111",
		230 => "01111111",
		231 => "01111111",
		232 => "01111111",
		233 => "01110010",
		234 => "11100000",
		235 => "01011111",
		236 => "01111111",
		237 => "01111111",
		238 => "01111111",
		239 => "01111111",
		240 => "01111111",
		241 => "01111011",
		242 => "11100000",
		243 => "01011111",
		244 => "01111111",
		245 => "01110011",
		246 => "11100000",
		247 => "01011010",
		248 => "11100000",
		249 => "01011010",
		250 => "11100000",
		251 => "11110000",


		-- Set the rest to zero
		others => x"00"
	);

begin

	q <= rom( to_integer( unsigned( addr ) ) );

end architecture;


--